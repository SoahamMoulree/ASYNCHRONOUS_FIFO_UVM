`define DSIZE 8
`define num_of_txns 100
`define ADDR 4
`define DEPTH 1 << 4
